// megafunction wizard: %FIR Compiler II v13.1%
// GENERATION: XML
// quad_bank_fir.v

// Generated using ACDS version 13.1 162 at 2015.02.20.23:46:16

`timescale 1 ps / 1 ps
module quad_bank_fir (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [13:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [34:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	quad_bank_fir_0002 quad_bank_fir_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2015 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="13.1" >
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone III" />
// Retrieval info: 	<generic name="filterType" value="Single Rate" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="L_bandsFilter" value="All taps" />
// Retrieval info: 	<generic name="clockRate" value="20" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="speedGrade" value="Medium" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="Read/Write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="symmetryMode" value="Symmetrical" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="inputRate" value=".08" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="inputType" value="Signed Binary" />
// Retrieval info: 	<generic name="inputBitWidth" value="12" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,-1.2251178286716597E-5,-9.155935311465223E-6,-1.2448394173141372E-5,-1.6419980964577204E-5,-2.1128353752928712E-5,-2.6634634507007285E-5,-3.3001642539319614E-5,-4.026804778490432E-5,-4.847865324283522E-5,-5.7651831772668165E-5,-6.780131943689444E-5,-7.892034819810176E-5,-9.098238073301963E-5,-1.0393522602367078E-4,-1.1770883087461122E-4,-1.3220306482073944E-4,-1.472907531296459E-4,-1.6281292688233857E-4,-1.7858082141795784E-4,-1.943727938349497E-4,-2.099362597736463E-4,-2.2498346537721384E-4,-2.3919578552993352E-4,-2.522230963875564E-4,-2.6368652050939585E-4,-2.73180031937078E-4,-2.802753580122796E-4,-2.8452319892380626E-4,-2.8545948922976223E-4,-2.8260985662295716E-4,-2.7549681360550666E-4,-2.6364567673750627E-4,-2.465921525177623E-4,-2.2388862610169194E-4,-1.9511406711927534E-4,-1.5988209544648646E-4,-1.1785051449988508E-4,-6.87301925021296E-5,-1.2294796436512277E-5,5.161103902559272E-5,1.230618820772515E-4,2.020432219680067E-4,2.88442580098405E-4,3.8204226968357205E-4,4.8251277840311133E-4,5.894077737376682E-4,7.021588526709495E-4,8.200727314410593E-4,9.423291308121401E-4,0.0010679806368393166,0.001195953994903435,0.0013250538478448482,0.0014539677400950506,0.0015812737337495618,0.001705449242003893,0.0018248823122275577,0.0019378848607132728,0.0020427080303572188,0.002137559035059679,0.002220620495761354,0.0022900710368865076,0.0023441074951612174,0.0023809681926005716,0.002398957407012291,0.002396470728421867,0.002372021356111042,0.002324266354949102,0.0022520331606769293,0.002154345717987916,0.002030449655007211,0.0018798363413768092,0.0017022657030062059,0.0014977872474357928,0.0012667590627699974,0.0010098642696478237,7.28124497244407E-4,4.229105764405792E-4,9.594962959077323E-5,-2.5067154389495647E-4,-6.145068354493161E-4,-9.927550891999245E-4,-0.0013822689930624377,-0.001779568063589901,-0.002180856390513248,-0.002582044347994294,-0.0029787746423283854,-0.003366452442179516,-0.0037402798572010805,-0.004095293573173398,-0.004426406816524127,-0.00472845415340425,-0.004996239277190043,-0.005224584771893611,-0.005408384349357559,-0.005542655951032734,-0.005622596692303996,-0.005643636953503348,-0.005601494570488072,-0.0054922278238397106,-0.005312287539578469,-0.005058566050683623,-0.004728445016338081,-0.00431983869473647,-0.003831233992264416,-0.0032617249666712306,-0.002611043048902999,-0.0018795807762438488,-0.001068411712409811,-1.7930185438096911E-4,7.852837130865266E-4,0.0018221815476998314,0.0029275365047565956,0.0040968178218316435,0.005324839671573426,0.006605791747514683,0.007933273587267474,0.00930033709768962,0.010699533131755295,0.012122966169324184,0.013562350790222123,0.015009080111994415,0.01645429337054208,0.01788894882117609,0.01930389552350913,0.020689952607576324,0.022037983133404895,0.023338979564043075,0.024584138721213743,0.02576494400291799,0.026873237718455005,0.027901297814453687,0.028841893373211684,0.02968837083934844,0.03043470645034635,0.031075568447292364,0.0316063430647714,0.03202321718142924,0.032323137022356535,0.032503981780977576,0.03256441750238264,0.032503981780977576,0.032323137022356535,0.03202321718142924,0.0316063430647714,0.031075568447292364,0.03043470645034635,0.02968837083934844,0.028841893373211684,0.027901297814453687,0.026873237718455005,0.02576494400291799,0.024584138721213743,0.023338979564043075,0.022037983133404895,0.020689952607576324,0.01930389552350913,0.01788894882117609,0.01645429337054208,0.015009080111994415,0.013562350790222123,0.012122966169324184,0.010699533131755295,0.00930033709768962,0.007933273587267474,0.006605791747514683,0.005324839671573426,0.0040968178218316435,0.0029275365047565956,0.0018221815476998314,7.852837130865266E-4,-1.7930185438096911E-4,-0.001068411712409811,-0.0018795807762438488,-0.002611043048902999,-0.0032617249666712306,-0.003831233992264416,-0.00431983869473647,-0.004728445016338081,-0.005058566050683623,-0.005312287539578469,-0.0054922278238397106,-0.005601494570488072,-0.005643636953503348,-0.005622596692303996,-0.005542655951032734,-0.005408384349357559,-0.005224584771893611,-0.004996239277190043,-0.00472845415340425,-0.004426406816524127,-0.004095293573173398,-0.0037402798572010805,-0.003366452442179516,-0.0029787746423283854,-0.002582044347994294,-0.002180856390513248,-0.001779568063589901,-0.0013822689930624377,-9.927550891999245E-4,-6.145068354493161E-4,-2.5067154389495647E-4,9.594962959077323E-5,4.229105764405792E-4,7.28124497244407E-4,0.0010098642696478237,0.0012667590627699974,0.0014977872474357928,0.0017022657030062059,0.0018798363413768092,0.002030449655007211,0.002154345717987916,0.0022520331606769293,0.002324266354949102,0.002372021356111042,0.002396470728421867,0.002398957407012291,0.0023809681926005716,0.0023441074951612174,0.0022900710368865076,0.002220620495761354,0.002137559035059679,0.0020427080303572188,0.0019378848607132728,0.0018248823122275577,0.001705449242003893,0.0015812737337495618,0.0014539677400950506,0.0013250538478448482,0.001195953994903435,0.0010679806368393166,9.423291308121401E-4,8.200727314410593E-4,7.021588526709495E-4,5.894077737376682E-4,4.8251277840311133E-4,3.8204226968357205E-4,2.88442580098405E-4,2.020432219680067E-4,1.230618820772515E-4,5.161103902559272E-5,-1.2294796436512277E-5,-6.87301925021296E-5,-1.1785051449988508E-4,-1.5988209544648646E-4,-1.9511406711927534E-4,-2.2388862610169194E-4,-2.465921525177623E-4,-2.6364567673750627E-4,-2.7549681360550666E-4,-2.8260985662295716E-4,-2.8545948922976223E-4,-2.8452319892380626E-4,-2.802753580122796E-4,-2.73180031937078E-4,-2.6368652050939585E-4,-2.522230963875564E-4,-2.3919578552993352E-4,-2.2498346537721384E-4,-2.099362597736463E-4,-1.943727938349497E-4,-1.7858082141795784E-4,-1.6281292688233857E-4,-1.472907531296459E-4,-1.3220306482073944E-4,-1.1770883087461122E-4,-1.0393522602367078E-4,-9.098238073301963E-5,-7.892034819810176E-5,-6.780131943689444E-5,-5.7651831772668165E-5,-4.847865324283522E-5,-4.026804778490432E-5,-3.3001642539319614E-5,-2.6634634507007285E-5,-2.1128353752928712E-5,-1.6419980964577204E-5,-1.2448394173141372E-5,-9.155935311465223E-6,-1.2251178286716597E-5,5.536261215769512E-4,3.990767727886767E-4,4.6863522455292206E-4,4.7895762697810313E-4,4.0555458198619093E-4,2.306269731523301E-4,-5.229625981724599E-5,-4.34202527594994E-4,-8.884073588572113E-4,-0.0013703651943626513,-0.0018204392726126422,-0.0021694630427440058,-0.002346681298486874,-0.0022896510156463017,-0.0019544677299845876,-0.0013251315328203191,-4.20536331786902E-4,7.02461734078238E-4,0.0019506016166222883,0.0032009510370268487,0.0043125758570195785,0.005142067642189852,0.005561278843086254,0.005475056454361597,0.004836548552886396,0.0036577487670162692,0.002013539887984898,3.807478211672226E-5,-0.0020867836838488287,-0.004149964220808589,-0.0059346557260363045,-0.007243942818502786,-0.00792538657874931,-0.00789129171234935,-0.007131716679921006,-0.005718062137164493,-0.0037962955121665417,-0.0015704643106065792,7.216307095535236E-4,0.00283766778952174,0.004561199195077909,0.00572903152360068,0.00625145050013258,0.006122676715051262,0.005420098045154586,0.004291731154822032,0.0029336136705462703,0.0015605925215860033,3.746985634547964E-4,-4.6495438484351974E-4,-8.657980446832519E-4,-8.145125206969183E-4,-3.7859021542769716E-4,3.049017047914505E-4,0.0010527976808250917,0.0016647346180574,0.0019579202985402504,0.0017978024999989715,0.001123121520031027,-4.045656409502689E-5,-0.0015804439389078668,-0.003310670408928678,-0.004997664049620507,-0.006394575606197093,-0.007279031693470181,-0.0074886319040237065,-0.0069479256082210575,-0.005683438787105456,-0.0038232491854595305,-0.0015807446583495804,7.749286165840522E-4,0.0029578701496096697,0.004708015333666661,0.0058305862819216635,0.006226076044072106,0.005905967272483812,0.004991222276995401,0.0036930979097047033,0.0022790981935269226,0.0010290640087343408,1.8802466098126515E-4,-7.658859756728052E-5,2.937817603701599E-4,0.0012345650903557513,0.0025637341039679573,0.004007358201485551,0.005241803244242087,0.005946412429926673,0.0058585604628612065,0.0048223046897448085,0.0028225273815891644,-1.7551202487881382E-6,-0.00336805386412358,-0.006884499867500726,-0.010103253122031615,-0.012585600420417386,-0.013968997854104973,-0.014025670432803141,-0.012703181598858995,-0.0101396111021489,-0.006649687616079597,-0.002683005726666643,0.001240712866338074,0.004610128991380656,0.007002486121378375,0.008153493877364073,0.008004731068021517,0.0067199782706728215,0.0046666642614331,0.0023625656965803018,3.951560489240541E-4,-6.756503244136912E-4,-4.183708442918468E-4,0.001386310752577628,0.004681957440558409,0.009122884178946399,0.014093596420193167,0.01878032837853721,0.022278344535023347,0.023720256541397047,0.022412752217224052,0.017960754003621873,0.01035848774369714,3.2661328491976206E-5,-0.012170574744263614,-0.025057029568351284,-0.03720913398951248,-0.04714981965151067,-0.05352545656713299,-0.055284430454171585,-0.05182760283923821,-0.04310998663793715,-0.029678173733429607,-0.012635937053296516,0.006460159520216277,0.02576407322214131,0.04334345062268734,0.05739820189258931,0.06646769412754208,0.06960084714332017,0.06646769412754208,0.05739820189258931,0.04334345062268734,0.02576407322214131,0.006460159520216277,-0.012635937053296516,-0.029678173733429607,-0.04310998663793715,-0.05182760283923821,-0.055284430454171585,-0.05352545656713299,-0.04714981965151067,-0.03720913398951248,-0.025057029568351284,-0.012170574744263614,3.2661328491976206E-5,0.01035848774369714,0.017960754003621873,0.022412752217224052,0.023720256541397047,0.022278344535023347,0.01878032837853721,0.014093596420193167,0.009122884178946399,0.004681957440558409,0.001386310752577628,-4.183708442918468E-4,-6.756503244136912E-4,3.951560489240541E-4,0.0023625656965803018,0.0046666642614331,0.0067199782706728215,0.008004731068021517,0.008153493877364073,0.007002486121378375,0.004610128991380656,0.001240712866338074,-0.002683005726666643,-0.006649687616079597,-0.0101396111021489,-0.012703181598858995,-0.014025670432803141,-0.013968997854104973,-0.012585600420417386,-0.010103253122031615,-0.006884499867500726,-0.00336805386412358,-1.7551202487881382E-6,0.0028225273815891644,0.0048223046897448085,0.0058585604628612065,0.005946412429926673,0.005241803244242087,0.004007358201485551,0.0025637341039679573,0.0012345650903557513,2.937817603701599E-4,-7.658859756728052E-5,1.8802466098126515E-4,0.0010290640087343408,0.0022790981935269226,0.0036930979097047033,0.004991222276995401,0.005905967272483812,0.006226076044072106,0.0058305862819216635,0.004708015333666661,0.0029578701496096697,7.749286165840522E-4,-0.0015807446583495804,-0.0038232491854595305,-0.005683438787105456,-0.0069479256082210575,-0.0074886319040237065,-0.007279031693470181,-0.006394575606197093,-0.004997664049620507,-0.003310670408928678,-0.0015804439389078668,-4.045656409502689E-5,0.001123121520031027,0.0017978024999989715,0.0019579202985402504,0.0016647346180574,0.0010527976808250917,3.049017047914505E-4,-3.7859021542769716E-4,-8.145125206969183E-4,-8.657980446832519E-4,-4.6495438484351974E-4,3.746985634547964E-4,0.0015605925215860033,0.0029336136705462703,0.004291731154822032,0.005420098045154586,0.006122676715051262,0.00625145050013258,0.00572903152360068,0.004561199195077909,0.00283766778952174,7.216307095535236E-4,-0.0015704643106065792,-0.0037962955121665417,-0.005718062137164493,-0.007131716679921006,-0.00789129171234935,-0.00792538657874931,-0.007243942818502786,-0.0059346557260363045,-0.004149964220808589,-0.0020867836838488287,3.807478211672226E-5,0.002013539887984898,0.0036577487670162692,0.004836548552886396,0.005475056454361597,0.005561278843086254,0.005142067642189852,0.0043125758570195785,0.0032009510370268487,0.0019506016166222883,7.02461734078238E-4,-4.20536331786902E-4,-0.0013251315328203191,-0.0019544677299845876,-0.0022896510156463017,-0.002346681298486874,-0.0021694630427440058,-0.0018204392726126422,-0.0013703651943626513,-8.884073588572113E-4,-4.34202527594994E-4,-5.229625981724599E-5,2.306269731523301E-4,4.0555458198619093E-4,4.7895762697810313E-4,4.6863522455292206E-4,3.990767727886767E-4,5.536261215769512E-4,0.011532487764135521,-0.05023338256322789,0.027647409743399107,0.02504331548917405,0.008846112413651097,-0.003779720504734646,-0.009982750400051924,-0.010870619923092687,-0.008390178292751417,-0.0043497573785606205,-1.5927756750550175E-4,0.0032166121594302596,0.005272970170183678,0.005901617612087814,0.005269046249962457,0.0037075077449052135,0.0016494159749679646,-4.6111031118168647E-4,-0.002268126047058724,-0.0035076245222607013,-0.004025487225961488,-0.0038297503265724083,-0.0030349943044470844,-0.0017996822560201458,-3.495891128884155E-4,0.001053492670510192,0.002211142314438503,0.00298136797979192,0.003255823465287068,0.0030305550019904897,0.0023640141549040403,0.0013476499701456604,1.68572563077159E-4,-0.0010021468490877905,-0.002018678284795935,-0.0027019991557336678,-0.0029908031287273758,-0.002841653023901497,-0.002254852084738464,-0.0013629763956393471,-2.5262739198318816E-4,8.697263316711266E-4,0.0018834394511034012,0.0026102202658484152,0.00296630645989003,0.002893104040644991,0.0024006611518928222,0.0015555317162308587,4.8098455292615837E-4,-6.795236609079392E-4,-0.0017569387353153561,-0.0026017605459449883,-0.003090207512487893,-0.0031381645292856246,-0.0027291976992785127,-0.001913602961878714,-8.008570911617227E-4,4.5638199675348753E-4,0.0016753357514791409,0.0026800338408742436,0.003325408286719878,0.0035001426765357757,0.0031691728854582137,0.0023719015908822373,0.001203341252914273,-1.731912843298789E-4,-0.001567398112616929,-0.0027837091031028753,-0.003632947619731863,-0.00398201507978696,-0.0037589105427487998,-0.0029720104394476607,-0.0017211254366259034,-1.724969692089358E-4,0.0014508818419520363,0.0029217331547433914,0.004014538972413889,0.004560292961212235,0.0044663341077720645,0.003717148367383366,0.0023901528993366897,6.615372030343381E-4,-0.0012486371623409364,-0.0030513393345799177,-0.004484744229396802,-0.005313254262193152,-0.005390521839787406,-0.00468239495751133,-0.003251759782817952,-0.0012886522536365652,9.579618947502162E-4,0.0031734906952855728,0.0050277395962096735,0.006244353019390433,0.006596797765342614,0.005984620612040909,0.0044590564121866514,0.0021874929068269526,-5.296874824877695E-4,-0.0033083470244594346,-0.0057521310274627,-0.007487082654314976,-0.008220728562669647,-0.007787166571968666,-0.006168671516770156,-0.003519575687560853,-1.7114906387460978E-4,0.003420378535743626,0.006745192116157484,0.009292239077966565,0.010640901451479848,0.010519095798961618,0.008817124111221741,0.005649407380075494,0.0013625986000724676,-0.0035008189426027144,-0.008284042588179948,-0.012238933494590081,-0.014764985061691823,-0.015259694131886502,-0.013617040248021309,-0.009575172778328278,-0.003712112004705064,0.0035741457705472184,0.011266500935909819,0.018262506941165248,0.023616175737259743,0.02616040299878552,0.0250306721774093,0.01976445953260703,0.010115168553594891,-0.0036331974710351084,-0.02065131949965968,-0.03988869781295981,-0.060045484822779535,-0.07948641827163644,-0.09655667935579067,-0.10990741854922989,-0.11846699214668578,0.8785734190893645,-0.11846699214668578,-0.10990741854922989,-0.09655667935579067,-0.07948641827163644,-0.060045484822779535,-0.03988869781295981,-0.02065131949965968,-0.0036331974710351084,0.010115168553594891,0.01976445953260703,0.0250306721774093,0.02616040299878552,0.023616175737259743,0.018262506941165248,0.011266500935909819,0.0035741457705472184,-0.003712112004705064,-0.009575172778328278,-0.013617040248021309,-0.015259694131886502,-0.014764985061691823,-0.012238933494590081,-0.008284042588179948,-0.0035008189426027144,0.0013625986000724676,0.005649407380075494,0.008817124111221741,0.010519095798961618,0.010640901451479848,0.009292239077966565,0.006745192116157484,0.003420378535743626,-1.7114906387460978E-4,-0.003519575687560853,-0.006168671516770156,-0.007787166571968666,-0.008220728562669647,-0.007487082654314976,-0.0057521310274627,-0.0033083470244594346,-5.296874824877695E-4,0.0021874929068269526,0.0044590564121866514,0.005984620612040909,0.006596797765342614,0.006244353019390433,0.0050277395962096735,0.0031734906952855728,9.579618947502162E-4,-0.0012886522536365652,-0.003251759782817952,-0.00468239495751133,-0.005390521839787406,-0.005313254262193152,-0.004484744229396802,-0.0030513393345799177,-0.0012486371623409364,6.615372030343381E-4,0.0023901528993366897,0.003717148367383366,0.0044663341077720645,0.004560292961212235,0.004014538972413889,0.0029217331547433914,0.0014508818419520363,-1.724969692089358E-4,-0.0017211254366259034,-0.0029720104394476607,-0.0037589105427487998,-0.00398201507978696,-0.003632947619731863,-0.0027837091031028753,-0.001567398112616929,-1.731912843298789E-4,0.001203341252914273,0.0023719015908822373,0.0031691728854582137,0.0035001426765357757,0.003325408286719878,0.0026800338408742436,0.0016753357514791409,4.5638199675348753E-4,-8.008570911617227E-4,-0.001913602961878714,-0.0027291976992785127,-0.0031381645292856246,-0.003090207512487893,-0.0026017605459449883,-0.0017569387353153561,-6.795236609079392E-4,4.8098455292615837E-4,0.0015555317162308587,0.0024006611518928222,0.002893104040644991,0.00296630645989003,0.0026102202658484152,0.0018834394511034012,8.697263316711266E-4,-2.5262739198318816E-4,-0.0013629763956393471,-0.002254852084738464,-0.002841653023901497,-0.0029908031287273758,-0.0027019991557336678,-0.002018678284795935,-0.0010021468490877905,1.68572563077159E-4,0.0013476499701456604,0.0023640141549040403,0.0030305550019904897,0.003255823465287068,0.00298136797979192,0.002211142314438503,0.001053492670510192,-3.495891128884155E-4,-0.0017996822560201458,-0.0030349943044470844,-0.0038297503265724083,-0.004025487225961488,-0.0035076245222607013,-0.002268126047058724,-4.6111031118168647E-4,0.0016494159749679646,0.0037075077449052135,0.005269046249962457,0.005901617612087814,0.005272970170183678,0.0032166121594302596,-1.5927756750550175E-4,-0.0043497573785606205,-0.008390178292751417,-0.010870619923092687,-0.009982750400051924,-0.003779720504734646,0.008846112413651097,0.02504331548917405,0.027647409743399107,-0.05023338256322789,0.011532487764135521" />
// Retrieval info: 	<generic name="coeffType" value="Signed Binary" />
// Retrieval info: 	<generic name="coeffScaling" value="Auto" />
// Retrieval info: 	<generic name="coeffBitWidth" value="14" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
// Retrieval info: 	<generic name="outType" value="Signed Binary" />
// Retrieval info: 	<generic name="outMSBRound" value="Saturating" />
// Retrieval info: 	<generic name="outMsbBitRem" value="0" />
// Retrieval info: 	<generic name="outLSBRound" value="Truncation" />
// Retrieval info: 	<generic name="outLsbBitRem" value="0" />
// Retrieval info: 	<generic name="resoureEstimation" value="1000,1200,10" />
// Retrieval info: 	<generic name="bankCount" value="4" />
// Retrieval info: 	<generic name="bankDisplay" value="3" />
// Retrieval info: </instance>
// IPFS_FILES : quad_bank_fir.vo
// RELATED_FILES: quad_bank_fir.v, altera_avalon_sc_fifo.v, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, dspba_library_package.vhd, dspba_library.vhd, quad_bank_fir_0002_rtl.vhd, quad_bank_fir_0002_ast.vhd, quad_bank_fir_0002.vhd
