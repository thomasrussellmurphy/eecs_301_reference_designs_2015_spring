//
// Copyright (c) 2015 Thomas R. Murphy and Case Western Reserve University
// All Rights Reserved
//
// Developed by Thomas Russell Murphy (trm70) during employment as teaching
// assistant of EECS 301 at CWRU.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS ``AS IS''
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR
// ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON
// ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//

module SEG7_LUT_4
       (
           input [ 15: 0 ] iDIG,
           output	[ 6: 0 ] oSEG0, oSEG1, oSEG2, oSEG3,
           output	oSEG0_DP, oSEG1_DP, oSEG2_DP, oSEG3_DP
       );


SEG7_LUT	u0	( oSEG0, oSEG0_DP, iDIG[ 3: 0 ] );
SEG7_LUT	u1	( oSEG1, oSEG1_DP, iDIG[ 7: 4 ] );
SEG7_LUT	u2	( oSEG2, oSEG2_DP, iDIG[ 11: 8 ] );
SEG7_LUT	u3	( oSEG3, oSEG3_DP, iDIG[ 15: 12 ] );

endmodule
