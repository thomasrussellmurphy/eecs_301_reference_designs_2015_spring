// megafunction wizard: %FIR Compiler II v13.1%
// GENERATION: XML
// quad_bank_fir.v

// Generated using ACDS version 13.1 162 at 2015.02.20.20:40:24

`timescale 1 ps / 1 ps
module quad_bank_fir (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [13:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [34:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	quad_bank_fir_0002 quad_bank_fir_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2015 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="13.1" >
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone III" />
// Retrieval info: 	<generic name="filterType" value="Single Rate" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="L_bandsFilter" value="All taps" />
// Retrieval info: 	<generic name="clockRate" value="20" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="speedGrade" value="Medium" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="Read/Write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="symmetryMode" value="Symmetrical" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="inputRate" value=".08" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="inputType" value="Signed Binary" />
// Retrieval info: 	<generic name="inputBitWidth" value="12" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,-1.2251178286716597E-5,-9.155935311465223E-6,-1.2448394173141372E-5,-1.6419980964577204E-5,-2.1128353752928712E-5,-2.6634634507007285E-5,-3.3001642539319614E-5,-4.026804778490432E-5,-4.847865324283522E-5,-5.7651831772668165E-5,-6.780131943689444E-5,-7.892034819810176E-5,-9.098238073301963E-5,-1.0393522602367078E-4,-1.1770883087461122E-4,-1.3220306482073944E-4,-1.472907531296459E-4,-1.6281292688233857E-4,-1.7858082141795784E-4,-1.943727938349497E-4,-2.099362597736463E-4,-2.2498346537721384E-4,-2.3919578552993352E-4,-2.522230963875564E-4,-2.6368652050939585E-4,-2.73180031937078E-4,-2.802753580122796E-4,-2.8452319892380626E-4,-2.8545948922976223E-4,-2.8260985662295716E-4,-2.7549681360550666E-4,-2.6364567673750627E-4,-2.465921525177623E-4,-2.2388862610169194E-4,-1.9511406711927534E-4,-1.5988209544648646E-4,-1.1785051449988508E-4,-6.87301925021296E-5,-1.2294796436512277E-5,5.161103902559272E-5,1.230618820772515E-4,2.020432219680067E-4,2.88442580098405E-4,3.8204226968357205E-4,4.8251277840311133E-4,5.894077737376682E-4,7.021588526709495E-4,8.200727314410593E-4,9.423291308121401E-4,0.0010679806368393166,0.001195953994903435,0.0013250538478448482,0.0014539677400950506,0.0015812737337495618,0.001705449242003893,0.0018248823122275577,0.0019378848607132728,0.0020427080303572188,0.002137559035059679,0.002220620495761354,0.0022900710368865076,0.0023441074951612174,0.0023809681926005716,0.002398957407012291,0.002396470728421867,0.002372021356111042,0.002324266354949102,0.0022520331606769293,0.002154345717987916,0.002030449655007211,0.0018798363413768092,0.0017022657030062059,0.0014977872474357928,0.0012667590627699974,0.0010098642696478237,7.28124497244407E-4,4.229105764405792E-4,9.594962959077323E-5,-2.5067154389495647E-4,-6.145068354493161E-4,-9.927550891999245E-4,-0.0013822689930624377,-0.001779568063589901,-0.002180856390513248,-0.002582044347994294,-0.0029787746423283854,-0.003366452442179516,-0.0037402798572010805,-0.004095293573173398,-0.004426406816524127,-0.00472845415340425,-0.004996239277190043,-0.005224584771893611,-0.005408384349357559,-0.005542655951032734,-0.005622596692303996,-0.005643636953503348,-0.005601494570488072,-0.0054922278238397106,-0.005312287539578469,-0.005058566050683623,-0.004728445016338081,-0.00431983869473647,-0.003831233992264416,-0.0032617249666712306,-0.002611043048902999,-0.0018795807762438488,-0.001068411712409811,-1.7930185438096911E-4,7.852837130865266E-4,0.0018221815476998314,0.0029275365047565956,0.0040968178218316435,0.005324839671573426,0.006605791747514683,0.007933273587267474,0.00930033709768962,0.010699533131755295,0.012122966169324184,0.013562350790222123,0.015009080111994415,0.01645429337054208,0.01788894882117609,0.01930389552350913,0.020689952607576324,0.022037983133404895,0.023338979564043075,0.024584138721213743,0.02576494400291799,0.026873237718455005,0.027901297814453687,0.028841893373211684,0.02968837083934844,0.03043470645034635,0.031075568447292364,0.0316063430647714,0.03202321718142924,0.032323137022356535,0.032503981780977576,0.03256441750238264,0.032503981780977576,0.032323137022356535,0.03202321718142924,0.0316063430647714,0.031075568447292364,0.03043470645034635,0.02968837083934844,0.028841893373211684,0.027901297814453687,0.026873237718455005,0.02576494400291799,0.024584138721213743,0.023338979564043075,0.022037983133404895,0.020689952607576324,0.01930389552350913,0.01788894882117609,0.01645429337054208,0.015009080111994415,0.013562350790222123,0.012122966169324184,0.010699533131755295,0.00930033709768962,0.007933273587267474,0.006605791747514683,0.005324839671573426,0.0040968178218316435,0.0029275365047565956,0.0018221815476998314,7.852837130865266E-4,-1.7930185438096911E-4,-0.001068411712409811,-0.0018795807762438488,-0.002611043048902999,-0.0032617249666712306,-0.003831233992264416,-0.00431983869473647,-0.004728445016338081,-0.005058566050683623,-0.005312287539578469,-0.0054922278238397106,-0.005601494570488072,-0.005643636953503348,-0.005622596692303996,-0.005542655951032734,-0.005408384349357559,-0.005224584771893611,-0.004996239277190043,-0.00472845415340425,-0.004426406816524127,-0.004095293573173398,-0.0037402798572010805,-0.003366452442179516,-0.0029787746423283854,-0.002582044347994294,-0.002180856390513248,-0.001779568063589901,-0.0013822689930624377,-9.927550891999245E-4,-6.145068354493161E-4,-2.5067154389495647E-4,9.594962959077323E-5,4.229105764405792E-4,7.28124497244407E-4,0.0010098642696478237,0.0012667590627699974,0.0014977872474357928,0.0017022657030062059,0.0018798363413768092,0.002030449655007211,0.002154345717987916,0.0022520331606769293,0.002324266354949102,0.002372021356111042,0.002396470728421867,0.002398957407012291,0.0023809681926005716,0.0023441074951612174,0.0022900710368865076,0.002220620495761354,0.002137559035059679,0.0020427080303572188,0.0019378848607132728,0.0018248823122275577,0.001705449242003893,0.0015812737337495618,0.0014539677400950506,0.0013250538478448482,0.001195953994903435,0.0010679806368393166,9.423291308121401E-4,8.200727314410593E-4,7.021588526709495E-4,5.894077737376682E-4,4.8251277840311133E-4,3.8204226968357205E-4,2.88442580098405E-4,2.020432219680067E-4,1.230618820772515E-4,5.161103902559272E-5,-1.2294796436512277E-5,-6.87301925021296E-5,-1.1785051449988508E-4,-1.5988209544648646E-4,-1.9511406711927534E-4,-2.2388862610169194E-4,-2.465921525177623E-4,-2.6364567673750627E-4,-2.7549681360550666E-4,-2.8260985662295716E-4,-2.8545948922976223E-4,-2.8452319892380626E-4,-2.802753580122796E-4,-2.73180031937078E-4,-2.6368652050939585E-4,-2.522230963875564E-4,-2.3919578552993352E-4,-2.2498346537721384E-4,-2.099362597736463E-4,-1.943727938349497E-4,-1.7858082141795784E-4,-1.6281292688233857E-4,-1.472907531296459E-4,-1.3220306482073944E-4,-1.1770883087461122E-4,-1.0393522602367078E-4,-9.098238073301963E-5,-7.892034819810176E-5,-6.780131943689444E-5,-5.7651831772668165E-5,-4.847865324283522E-5,-4.026804778490432E-5,-3.3001642539319614E-5,-2.6634634507007285E-5,-2.1128353752928712E-5,-1.6419980964577204E-5,-1.2448394173141372E-5,-9.155935311465223E-6,-1.2251178286716597E-5,5.536261215769512E-4,3.990767727886767E-4,4.6863522455292206E-4,4.7895762697810313E-4,4.0555458198619093E-4,2.306269731523301E-4,-5.229625981724599E-5,-4.34202527594994E-4,-8.884073588572113E-4,-0.0013703651943626513,-0.0018204392726126422,-0.0021694630427440058,-0.002346681298486874,-0.0022896510156463017,-0.0019544677299845876,-0.0013251315328203191,-4.20536331786902E-4,7.02461734078238E-4,0.0019506016166222883,0.0032009510370268487,0.0043125758570195785,0.005142067642189852,0.005561278843086254,0.005475056454361597,0.004836548552886396,0.0036577487670162692,0.002013539887984898,3.807478211672226E-5,-0.0020867836838488287,-0.004149964220808589,-0.0059346557260363045,-0.007243942818502786,-0.00792538657874931,-0.00789129171234935,-0.007131716679921006,-0.005718062137164493,-0.0037962955121665417,-0.0015704643106065792,7.216307095535236E-4,0.00283766778952174,0.004561199195077909,0.00572903152360068,0.00625145050013258,0.006122676715051262,0.005420098045154586,0.004291731154822032,0.0029336136705462703,0.0015605925215860033,3.746985634547964E-4,-4.6495438484351974E-4,-8.657980446832519E-4,-8.145125206969183E-4,-3.7859021542769716E-4,3.049017047914505E-4,0.0010527976808250917,0.0016647346180574,0.0019579202985402504,0.0017978024999989715,0.001123121520031027,-4.045656409502689E-5,-0.0015804439389078668,-0.003310670408928678,-0.004997664049620507,-0.006394575606197093,-0.007279031693470181,-0.0074886319040237065,-0.0069479256082210575,-0.005683438787105456,-0.0038232491854595305,-0.0015807446583495804,7.749286165840522E-4,0.0029578701496096697,0.004708015333666661,0.0058305862819216635,0.006226076044072106,0.005905967272483812,0.004991222276995401,0.0036930979097047033,0.0022790981935269226,0.0010290640087343408,1.8802466098126515E-4,-7.658859756728052E-5,2.937817603701599E-4,0.0012345650903557513,0.0025637341039679573,0.004007358201485551,0.005241803244242087,0.005946412429926673,0.0058585604628612065,0.0048223046897448085,0.0028225273815891644,-1.7551202487881382E-6,-0.00336805386412358,-0.006884499867500726,-0.010103253122031615,-0.012585600420417386,-0.013968997854104973,-0.014025670432803141,-0.012703181598858995,-0.0101396111021489,-0.006649687616079597,-0.002683005726666643,0.001240712866338074,0.004610128991380656,0.007002486121378375,0.008153493877364073,0.008004731068021517,0.0067199782706728215,0.0046666642614331,0.0023625656965803018,3.951560489240541E-4,-6.756503244136912E-4,-4.183708442918468E-4,0.001386310752577628,0.004681957440558409,0.009122884178946399,0.014093596420193167,0.01878032837853721,0.022278344535023347,0.023720256541397047,0.022412752217224052,0.017960754003621873,0.01035848774369714,3.2661328491976206E-5,-0.012170574744263614,-0.025057029568351284,-0.03720913398951248,-0.04714981965151067,-0.05352545656713299,-0.055284430454171585,-0.05182760283923821,-0.04310998663793715,-0.029678173733429607,-0.012635937053296516,0.006460159520216277,0.02576407322214131,0.04334345062268734,0.05739820189258931,0.06646769412754208,0.06960084714332017,0.06646769412754208,0.05739820189258931,0.04334345062268734,0.02576407322214131,0.006460159520216277,-0.012635937053296516,-0.029678173733429607,-0.04310998663793715,-0.05182760283923821,-0.055284430454171585,-0.05352545656713299,-0.04714981965151067,-0.03720913398951248,-0.025057029568351284,-0.012170574744263614,3.2661328491976206E-5,0.01035848774369714,0.017960754003621873,0.022412752217224052,0.023720256541397047,0.022278344535023347,0.01878032837853721,0.014093596420193167,0.009122884178946399,0.004681957440558409,0.001386310752577628,-4.183708442918468E-4,-6.756503244136912E-4,3.951560489240541E-4,0.0023625656965803018,0.0046666642614331,0.0067199782706728215,0.008004731068021517,0.008153493877364073,0.007002486121378375,0.004610128991380656,0.001240712866338074,-0.002683005726666643,-0.006649687616079597,-0.0101396111021489,-0.012703181598858995,-0.014025670432803141,-0.013968997854104973,-0.012585600420417386,-0.010103253122031615,-0.006884499867500726,-0.00336805386412358,-1.7551202487881382E-6,0.0028225273815891644,0.0048223046897448085,0.0058585604628612065,0.005946412429926673,0.005241803244242087,0.004007358201485551,0.0025637341039679573,0.0012345650903557513,2.937817603701599E-4,-7.658859756728052E-5,1.8802466098126515E-4,0.0010290640087343408,0.0022790981935269226,0.0036930979097047033,0.004991222276995401,0.005905967272483812,0.006226076044072106,0.0058305862819216635,0.004708015333666661,0.0029578701496096697,7.749286165840522E-4,-0.0015807446583495804,-0.0038232491854595305,-0.005683438787105456,-0.0069479256082210575,-0.0074886319040237065,-0.007279031693470181,-0.006394575606197093,-0.004997664049620507,-0.003310670408928678,-0.0015804439389078668,-4.045656409502689E-5,0.001123121520031027,0.0017978024999989715,0.0019579202985402504,0.0016647346180574,0.0010527976808250917,3.049017047914505E-4,-3.7859021542769716E-4,-8.145125206969183E-4,-8.657980446832519E-4,-4.6495438484351974E-4,3.746985634547964E-4,0.0015605925215860033,0.0029336136705462703,0.004291731154822032,0.005420098045154586,0.006122676715051262,0.00625145050013258,0.00572903152360068,0.004561199195077909,0.00283766778952174,7.216307095535236E-4,-0.0015704643106065792,-0.0037962955121665417,-0.005718062137164493,-0.007131716679921006,-0.00789129171234935,-0.00792538657874931,-0.007243942818502786,-0.0059346557260363045,-0.004149964220808589,-0.0020867836838488287,3.807478211672226E-5,0.002013539887984898,0.0036577487670162692,0.004836548552886396,0.005475056454361597,0.005561278843086254,0.005142067642189852,0.0043125758570195785,0.0032009510370268487,0.0019506016166222883,7.02461734078238E-4,-4.20536331786902E-4,-0.0013251315328203191,-0.0019544677299845876,-0.0022896510156463017,-0.002346681298486874,-0.0021694630427440058,-0.0018204392726126422,-0.0013703651943626513,-8.884073588572113E-4,-4.34202527594994E-4,-5.229625981724599E-5,2.306269731523301E-4,4.0555458198619093E-4,4.7895762697810313E-4,4.6863522455292206E-4,3.990767727886767E-4,5.536261215769512E-4,8.99204136193031E-4,-0.0029575027410878607,0.0012522259330968518,0.0014474715355132352,6.153603854221618E-4,-1.659931881556894E-4,-5.986731256551441E-4,-6.863956045071775E-4,-5.311108928363826E-4,-2.511867672212154E-4,5.1324131103023544E-5,3.007637811312996E-4,4.495736657970332E-4,4.775407744281502E-4,3.894993578087353E-4,2.1098059398066832E-4,-1.6312490029624014E-5,-2.4096305333386146E-4,-4.131163526204453E-4,-4.925854121350706E-4,-4.568968066005983E-4,-3.099440830397532E-4,-8.040061542205302E-5,1.827968352032964E-4,4.179583360227206E-4,5.667486955231765E-4,5.871568227751245E-4,4.6497624376681205E-4,2.209490675408872E-4,-9.491383734098202E-5,-4.1065312536942586E-4,-6.485535418477783E-4,-7.456740879833271E-4,-6.669132967575787E-4,-4.2000264986531786E-4,-5.0839905098100464E-5,3.5793402378033693E-4,7.100758113420829E-4,9.140190264703736E-4,9.096405677768592E-4,6.824017941375739E-4,2.726514286011081E-4,-2.3320723769062118E-4,-7.181701121643318E-4,-0.0010631981291398145,-0.0011751302495203856,-0.0010101687494916026,-5.889090233827862E-4,5.1105012068968994E-6,6.40026322219895E-4,0.00116424702232121,0.0014429831172431105,0.0013920919855901304,0.0010022421085057946,3.447891711178826E-4,-4.402712331484532E-4,-0.0011725060046616903,-0.0016724867911583085,-0.0018041536996896777,-0.0015108801391846437,-8.353602653674448E-4,8.526515913275322E-5,0.0010453122112885785,0.0018170663930551524,0.0022048679887921845,0.002091198247725927,0.00147064886667169,4.577038432151147E-4,-7.298545296808244E-4,-0.0018196375304654873,-0.002543116593769817,-0.0027077523447254464,-0.002237195843737918,-0.0012063133947472267,1.793404612346655E-4,0.0016098735655041745,0.002748196421947866,0.0033045240956368323,0.00310994694850826,0.0021666751610468155,6.48818634490311E-4,-0.001121260997070998,-0.0027366854073748287,-0.003804290310178759,-0.004037302823850845,-0.0033288584407518778,-0.0017867483442603573,2.798505279261117E-4,0.002413686813651156,0.00411079069931715,0.00494473446073284,0.004664345555261978,0.003258418527894764,9.855527772395774E-4,-0.001668616084221464,-0.004105558050679065,-0.005738386582495487,-0.00611984319607265,-0.005076487074326291,-0.0027619087319974223,3.747311435897348E-4,0.0036461816529379126,0.006284942902895052,0.007633069652197109,0.0072619809264840825,0.005145848160771344,0.0016398722791234805,-0.0025279702357895863,-0.006429082969330111,-0.009117507936553717,-0.009859689083604876,-0.008315258186701636,-0.004651447512844679,4.528883874126907E-4,0.005920871066257214,0.010493476525566073,0.013002089162310243,0.012645545091794936,0.009210003312702688,0.0031756985946148767,-0.004320025844066372,-0.011672835058134162,-0.017123046016091617,-0.019130728517354416,-0.016746296230240387,-0.009893102390777815,5.03547533176785E-4,0.012577827071151427,0.023782861056838307,0.03130845752243827,0.0325889677096637,0.02581124584465437,0.010321502545721947,-0.013147591845476727,-0.04248564398210944,-0.07445720178938144,-0.10516073570420158,-0.13062769723541479,-0.14744782316317936,0.8466752209601254,-0.14744782316317936,-0.13062769723541479,-0.10516073570420158,-0.07445720178938144,-0.04248564398210944,-0.013147591845476727,0.010321502545721947,0.02581124584465437,0.0325889677096637,0.03130845752243827,0.023782861056838307,0.012577827071151427,5.03547533176785E-4,-0.009893102390777815,-0.016746296230240387,-0.019130728517354416,-0.017123046016091617,-0.011672835058134162,-0.004320025844066372,0.0031756985946148767,0.009210003312702688,0.012645545091794936,0.013002089162310243,0.010493476525566073,0.005920871066257214,4.528883874126907E-4,-0.004651447512844679,-0.008315258186701636,-0.009859689083604876,-0.009117507936553717,-0.006429082969330111,-0.0025279702357895863,0.0016398722791234805,0.005145848160771344,0.0072619809264840825,0.007633069652197109,0.006284942902895052,0.0036461816529379126,3.747311435897348E-4,-0.0027619087319974223,-0.005076487074326291,-0.00611984319607265,-0.005738386582495487,-0.004105558050679065,-0.001668616084221464,9.855527772395774E-4,0.003258418527894764,0.004664345555261978,0.00494473446073284,0.00411079069931715,0.002413686813651156,2.798505279261117E-4,-0.0017867483442603573,-0.0033288584407518778,-0.004037302823850845,-0.003804290310178759,-0.0027366854073748287,-0.001121260997070998,6.48818634490311E-4,0.0021666751610468155,0.00310994694850826,0.0033045240956368323,0.002748196421947866,0.0016098735655041745,1.793404612346655E-4,-0.0012063133947472267,-0.002237195843737918,-0.0027077523447254464,-0.002543116593769817,-0.0018196375304654873,-7.298545296808244E-4,4.577038432151147E-4,0.00147064886667169,0.002091198247725927,0.0022048679887921845,0.0018170663930551524,0.0010453122112885785,8.526515913275322E-5,-8.353602653674448E-4,-0.0015108801391846437,-0.0018041536996896777,-0.0016724867911583085,-0.0011725060046616903,-4.402712331484532E-4,3.447891711178826E-4,0.0010022421085057946,0.0013920919855901304,0.0014429831172431105,0.00116424702232121,6.40026322219895E-4,5.1105012068968994E-6,-5.889090233827862E-4,-0.0010101687494916026,-0.0011751302495203856,-0.0010631981291398145,-7.181701121643318E-4,-2.3320723769062118E-4,2.726514286011081E-4,6.824017941375739E-4,9.096405677768592E-4,9.140190264703736E-4,7.100758113420829E-4,3.5793402378033693E-4,-5.0839905098100464E-5,-4.2000264986531786E-4,-6.669132967575787E-4,-7.456740879833271E-4,-6.485535418477783E-4,-4.1065312536942586E-4,-9.491383734098202E-5,2.209490675408872E-4,4.6497624376681205E-4,5.871568227751245E-4,5.667486955231765E-4,4.179583360227206E-4,1.827968352032964E-4,-8.040061542205302E-5,-3.099440830397532E-4,-4.568968066005983E-4,-4.925854121350706E-4,-4.131163526204453E-4,-2.4096305333386146E-4,-1.6312490029624014E-5,2.1098059398066832E-4,3.894993578087353E-4,4.775407744281502E-4,4.495736657970332E-4,3.007637811312996E-4,5.1324131103023544E-5,-2.511867672212154E-4,-5.311108928363826E-4,-6.863956045071775E-4,-5.986731256551441E-4,-1.659931881556894E-4,6.153603854221618E-4,0.0014474715355132352,0.0012522259330968518,-0.0029575027410878607,8.99204136193031E-4" />
// Retrieval info: 	<generic name="coeffType" value="Signed Binary" />
// Retrieval info: 	<generic name="coeffScaling" value="Auto" />
// Retrieval info: 	<generic name="coeffBitWidth" value="14" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
// Retrieval info: 	<generic name="outType" value="Signed Binary" />
// Retrieval info: 	<generic name="outMSBRound" value="Saturating" />
// Retrieval info: 	<generic name="outMsbBitRem" value="0" />
// Retrieval info: 	<generic name="outLSBRound" value="Truncation" />
// Retrieval info: 	<generic name="outLsbBitRem" value="0" />
// Retrieval info: 	<generic name="resoureEstimation" value="1000,1200,10" />
// Retrieval info: 	<generic name="bankCount" value="4" />
// Retrieval info: 	<generic name="bankDisplay" value="3" />
// Retrieval info: </instance>
// IPFS_FILES : quad_bank_fir.vo
// RELATED_FILES: quad_bank_fir.v, altera_avalon_sc_fifo.v, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, dspba_library_package.vhd, dspba_library.vhd, quad_bank_fir_0002_rtl.vhd, quad_bank_fir_0002_ast.vhd, quad_bank_fir_0002.vhd
