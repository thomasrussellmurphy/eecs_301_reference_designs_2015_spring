// megafunction wizard: %FIR Compiler II v13.1%
// GENERATION: XML
// fir_hpf.v

// Generated using ACDS version 13.1 162 at 2015.04.14.23:27:54

`timescale 1 ps / 1 ps
module fir_hpf (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [11:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [11:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	fir_hpf_0002 fir_hpf_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2015 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="13.1" >
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone III" />
// Retrieval info: 	<generic name="filterType" value="Single Rate" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="L_bandsFilter" value="All taps" />
// Retrieval info: 	<generic name="clockRate" value="50" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="speedGrade" value="Medium" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="Read/Write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="symmetryMode" value="Non Symmetry" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="inputRate" value=".05" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="inputType" value="Signed Binary" />
// Retrieval info: 	<generic name="inputBitWidth" value="12" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="0.0,0.0,0.0,0.0,0.0,1.28746E-6,1.82361E-6,2.43071E-6,3.09494E-6,3.79927E-6,4.52541E-6,5.25146E-6,5.95503E-6,6.60968E-6,7.18944E-6,7.66376E-6,8.00378E-6,8.1755E-6,8.14804E-6,7.88473E-6,7.35374E-6,6.5167E-6,5.34206E-6,3.79093E-6,1.83343E-6,0.0,-3.44153E-6,-6.8214E-6,-1.07298E-5,-1.51986E-5,-2.02426E-5,-2.58881E-5,-3.21412E-5,-3.90209E-5,-4.65225E-5,-5.46558E-5,-6.34036E-5,-7.27648E-5,-8.27077E-5,-9.32188E-5,-1.0425E-4,-1.15774E-4,-1.27726E-4,-1.40063E-4,-1.527E-4,-1.65581E-4,-1.786E-4,-1.91684E-4,-2.04708E-4,-2.17584E-4,-2.30167E-4,-2.42354E-4,-2.5398E-4,-2.64928E-4,-2.75018E-4,-2.84121E-4,-2.92041E-4,-2.98641E-4,-3.03712E-4,-3.07112E-4,-3.08625E-4,-3.08108E-4,-3.05339E-4,-3.00181E-4,-2.92414E-4,-2.81909E-4,-2.68452E-4,-2.51933E-4,-2.32151E-4,-2.09016E-4,-1.82346E-4,-1.52085E-4,-1.18075E-4,-8.02948E-5,-3.86222E-5,6.92031E-6,5.64161E-5,1.09791E-4,1.67084E-4,2.28161E-4,2.9301E-4,3.61436E-4,4.33368E-4,5.08542E-4,5.86828E-4,6.6789E-4,7.51533E-4,8.37347E-4,9.25071E-4,0.00101422,0.00110447,0.00119526,0.0012862,0.00137665,0.00146618,0.00155407,0.00163982,0.00172267,0.00180206,0.00187718,0.00194744,0.00201197,0.00207016,0.00212111,0.00216418,0.00219847,0.00222332,0.00223784,0.00224138,0.00223304,0.00221224,0.00217808,0.00213002,0.00206722,0.00198919,0.00189517,0.00178475,0.00165722,0.00151229,0.00134935,0.0011682,9.68354E-4,7.49744E-4,5.11994E-4,2.55185E-4,-2.09265E-5,-3.1611E-4,-6.30461E-4,-9.63593E-4,-0.00131545,-0.00168548,-0.00207346,-0.00247869,-0.00290079,-0.00333887,-0.00379241,-0.00426036,-0.00474204,-0.00523624,-0.00574215,-0.00625842,-0.0067841,-0.0073177,-0.00785816,-0.00840388,-0.00895369,-0.0095059,-0.0100593,-0.010612,-0.0111629,-0.01171,-0.012252,-0.0127871,-0.013314,-0.0138307,-0.014336,-0.0148281,-0.0153057,-0.015767,-0.0162108,-0.0166354,-0.0170397,-0.0174222,-0.0177818,-0.0181172,-0.0184274,-0.0187111,-0.0189678,-0.0191962,-0.0193959,-0.0195658,-0.0197058,-0.0198151,-0.0198935,-0.0199406,0.979323,-0.0199406,-0.0198935,-0.0198151,-0.0197058,-0.0195658,-0.0193959,-0.0191962,-0.0189678,-0.0187111,-0.0184274,-0.0181172,-0.0177818,-0.0174222,-0.0170397,-0.0166354,-0.0162108,-0.015767,-0.0153057,-0.0148281,-0.014336,-0.0138307,-0.013314,-0.0127871,-0.012252,-0.01171,-0.0111629,-0.010612,-0.0100593,-0.0095059,-0.00895369,-0.00840388,-0.00785816,-0.0073177,-0.0067841,-0.00625842,-0.00574215,-0.00523624,-0.00474204,-0.00426036,-0.00379241,-0.00333887,-0.00290079,-0.00247869,-0.00207346,-0.00168548,-0.00131545,-9.63593E-4,-6.30461E-4,-3.1611E-4,-2.09265E-5,2.55185E-4,5.11994E-4,7.49744E-4,9.68354E-4,0.0011682,0.00134935,0.00151229,0.00165722,0.00178475,0.00189517,0.00198919,0.00206722,0.00213002,0.00217808,0.00221224,0.00223304,0.00224138,0.00223784,0.00222332,0.00219847,0.00216418,0.00212111,0.00207016,0.00201197,0.00194744,0.00187718,0.00180206,0.00172267,0.00163982,0.00155407,0.00146618,0.00137665,0.0012862,0.00119526,0.00110447,0.00101422,9.25071E-4,8.37347E-4,7.51533E-4,6.6789E-4,5.86828E-4,5.08542E-4,4.33368E-4,3.61436E-4,2.9301E-4,2.28161E-4,1.67084E-4,1.09791E-4,5.64161E-5,6.92031E-6,-3.86222E-5,-8.02948E-5,-1.18075E-4,-1.52085E-4,-1.82346E-4,-2.09016E-4,-2.32151E-4,-2.51933E-4,-2.68452E-4,-2.81909E-4,-2.92414E-4,-3.00181E-4,-3.05339E-4,-3.08108E-4,-3.08625E-4,-3.07112E-4,-3.03712E-4,-2.98641E-4,-2.92041E-4,-2.84121E-4,-2.75018E-4,-2.64928E-4,-2.5398E-4,-2.42354E-4,-2.30167E-4,-2.17584E-4,-2.04708E-4,-1.91684E-4,-1.786E-4,-1.65581E-4,-1.527E-4,-1.40063E-4,-1.27726E-4,-1.15774E-4,-1.0425E-4,-9.32188E-5,-8.27077E-5,-7.27648E-5,-6.34036E-5,-5.46558E-5,-4.65225E-5,-3.90209E-5,-3.21412E-5,-2.58881E-5,-2.02426E-5,-1.51986E-5,-1.07298E-5,-6.8214E-6,-3.44153E-6,0.0,1.83343E-6,3.79093E-6,5.34206E-6,6.5167E-6,7.35374E-6,7.88473E-6,8.14804E-6,8.1755E-6,8.00378E-6,7.66376E-6,7.18944E-6,6.60968E-6,5.95503E-6,5.25146E-6,4.52541E-6,3.79927E-6,3.09494E-6,2.43071E-6,1.82361E-6,1.28746E-6,0.0,0.0,0.0,0.0,0.0" />
// Retrieval info: 	<generic name="coeffType" value="Signed Binary" />
// Retrieval info: 	<generic name="coeffScaling" value="Auto" />
// Retrieval info: 	<generic name="coeffBitWidth" value="16" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
// Retrieval info: 	<generic name="outType" value="Signed Binary" />
// Retrieval info: 	<generic name="outMSBRound" value="Saturating" />
// Retrieval info: 	<generic name="outMsbBitRem" value="9" />
// Retrieval info: 	<generic name="outLSBRound" value="Truncation" />
// Retrieval info: 	<generic name="outLsbBitRem" value="16" />
// Retrieval info: 	<generic name="resoureEstimation" value="1000,1200,10" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : fir_hpf.vo
// RELATED_FILES: fir_hpf.v, altera_avalon_sc_fifo.v, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, dspba_library_package.vhd, dspba_library.vhd, fir_hpf_0002_rtl.vhd, fir_hpf_0002_ast.vhd, fir_hpf_0002.vhd
