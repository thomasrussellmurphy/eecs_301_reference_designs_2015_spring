// megafunction wizard: %FIR Compiler II v13.1%
// GENERATION: XML
// fir_lpf.v

// Generated using ACDS version 13.1 162 at 2015.04.15.13:22:42

`timescale 1 ps / 1 ps
module fir_lpf (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [11:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [11:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	fir_lpf_0002 fir_lpf_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2015 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="13.1" >
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone III" />
// Retrieval info: 	<generic name="filterType" value="Single Rate" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="L_bandsFilter" value="All taps" />
// Retrieval info: 	<generic name="clockRate" value="20" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="speedGrade" value="Medium" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="Read/Write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="symmetryMode" value="Non Symmetry" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="inputRate" value=".05" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="inputType" value="Signed Binary" />
// Retrieval info: 	<generic name="inputBitWidth" value="12" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="-9.314227689476197E-5,-8.791028569757087E-6,-8.607316290639185E-6,-7.973763240331752E-6,-6.843685137216114E-6,-5.1627963389752305E-6,-2.8782725794033763E-6,6.773457347335861E-8,3.7340395101024115E-6,8.181670695133963E-6,1.3474034479830275E-5,1.967652583693631E-5,2.685486721875701E-5,3.5075205134138346E-5,4.440230106207581E-5,5.489773300334159E-5,6.662077754901276E-5,7.962974039102439E-5,9.398288772764757E-5,1.0973572173158561E-4,1.2693578037493446E-4,1.4561660801765025E-4,1.6580895365819176E-4,1.8755202781569998E-4,2.108893983098659E-4,2.3578135519507906E-4,2.6228274935093744E-4,2.903616395363066E-4,3.200137461957706E-4,3.5120864671016344E-4,3.8391283512202143E-4,4.180750727639507E-4,4.536340834518712E-4,4.905157202469902E-4,5.286317701011066E-4,5.678804755293912E-4,6.081483601883429E-4,6.493072085284562E-4,6.912130516169605E-4,7.337077975763362E-4,7.766209124107469E-4,8.197694451210797E-4,8.62955798960464E-4,9.059666182415098E-4,9.485751242191463E-4,9.905471698109832E-4,0.0010316369578531872,0.0010715828256110285,0.0011101104561474747,0.00114695406560225,0.001181814956554507,0.0012144105515198558,0.0012444355144887226,0.0012715955672936968,0.0012955794786071852,0.0013160876400487337,0.0013328148472630697,0.0013454577372516694,0.0013537200572276192,0.0013573134214608581,0.001355954523788637,0.0013493699157382595,0.0013373001969577845,0.0013195016209159504,0.0012957461488201504,0.0012658227447402998,0.0012295408339795142,0.0011867342580300108,0.0011372628442138308,0.0010810102355067698,0.0010178880877549088,9.478404676130159E-4,8.70844964072757E-4,7.86906446323214E-4,6.960756385164889E-4,5.984277236095604E-4,4.940920673403825E-4,3.8321319301009194E-4,2.6601121168961974E-4,1.4271233464115002E-4,1.3603335227636716E-5,-1.2098390162180816E-4,-2.606803675417535E-4,-4.050781679815073E-4,-5.537220980725372E-4,-7.06112330338158E-4,-8.617084696593745E-4,-0.00101993169925511,-0.0011801639173750279,-0.0013417471650933996,-0.0015039847400529322,-0.001666144828375941,-0.0018274637060259303,-0.0019871455436864063,-0.0021443652375523884,-0.0022982715177295777,-0.0024479897165633497,-0.002592621567003264,-0.0027312567521084546,-0.002862962330892213,-0.002986827340128685,-0.003101831706927529,-0.003207161130732031,-0.0033017673961671288,-0.0033847288158777504,-0.0034551415290471933,-0.003512100725539874,-0.0035547056081431157,-0.0035820790299364172,-0.00359337524746581,-0.003587784109429537,-0.003564532401333533,-0.0035228861172754804,-0.0034621539402339366,-0.0033816936183415428,-0.0032809176021118686,-0.0031592976392567315,-0.0030163699464840297,-0.002851737169858066,-0.002665068345937549,-0.002456096750531026,-0.002224619181984385,-0.001970493049077555,-0.0016936559390717152,-0.0013941676049199915,-0.001072456045279717,-7.28185739138134E-4,-3.6203177202829797E-4,2.5743555612137195E-5,4.3466095821653386E-4,8.641708058785863E-4,0.0013136341318983284,0.0017823306649008331,0.0022694557392816156,0.0027741222712723583,0.0032953631556954504,0.0038321339979232975,0.004383314684813668,0.004947714248015303,0.005524074381750709,0.006111070991248544,0.006707317032396235,0.007311367429232032,0.007921727018075494,0.008536857528040242,0.009155180777909258,0.009775074467086697,0.010394882233693628,0.011012932189119267,0.01162755209127645,0.01223700491497296,0.012839606531884297,0.013433631708801833,0.014017383965648797,0.014589167194400694,0.015147314371887065,0.01569017826261504,0.016216146378403396,0.016723645877498618,0.017211147668940125,0.01767717233992148,0.018120299891767156,0.018539173805098497,0.01893250426131548,0.019299073349307413,0.01963774177286249,0.01994745492859834,0.020227245905441307,0.02047623678985522,0.020693641615178875,0.020878775698108892,0.02103105693236326,0.021150003025647547,0.02123523114835423,0.02128648059189456,0.021303579101765974,0.02128648059189456,0.02123523114835423,0.021150003025647547,0.02103105693236326,0.020878775698108892,0.020693641615178875,0.02047623678985522,0.020227245905441307,0.01994745492859834,0.01963774177286249,0.019299073349307413,0.01893250426131548,0.018539173805098497,0.018120299891767156,0.01767717233992148,0.017211147668940125,0.016723645877498618,0.016216146378403396,0.01569017826261504,0.015147314371887065,0.014589167194400694,0.014017383965648797,0.013433631708801833,0.012839606531884297,0.01223700491497296,0.01162755209127645,0.011012932189119267,0.010394882233693628,0.009775074467086697,0.009155180777909258,0.008536857528040242,0.007921727018075494,0.007311367429232032,0.006707317032396235,0.006111070991248544,0.005524074381750709,0.004947714248015303,0.004383314684813668,0.0038321339979232975,0.0032953631556954504,0.0027741222712723583,0.0022694557392816156,0.0017823306649008331,0.0013136341318983284,8.641708058785863E-4,4.3466095821653386E-4,2.5743555612137195E-5,-3.6203177202829797E-4,-7.28185739138134E-4,-0.001072456045279717,-0.0013941676049199915,-0.0016936559390717152,-0.001970493049077555,-0.002224619181984385,-0.002456096750531026,-0.002665068345937549,-0.002851737169858066,-0.0030163699464840297,-0.0031592976392567315,-0.0032809176021118686,-0.0033816936183415428,-0.0034621539402339366,-0.0035228861172754804,-0.003564532401333533,-0.003587784109429537,-0.00359337524746581,-0.0035820790299364172,-0.0035547056081431157,-0.003512100725539874,-0.0034551415290471933,-0.0033847288158777504,-0.0033017673961671288,-0.003207161130732031,-0.003101831706927529,-0.002986827340128685,-0.002862962330892213,-0.0027312567521084546,-0.002592621567003264,-0.0024479897165633497,-0.0022982715177295777,-0.0021443652375523884,-0.0019871455436864063,-0.0018274637060259303,-0.001666144828375941,-0.0015039847400529322,-0.0013417471650933996,-0.0011801639173750279,-0.00101993169925511,-8.617084696593745E-4,-7.06112330338158E-4,-5.537220980725372E-4,-4.050781679815073E-4,-2.606803675417535E-4,-1.2098390162180816E-4,1.3603335227636716E-5,1.4271233464115002E-4,2.6601121168961974E-4,3.8321319301009194E-4,4.940920673403825E-4,5.984277236095604E-4,6.960756385164889E-4,7.86906446323214E-4,8.70844964072757E-4,9.478404676130159E-4,0.0010178880877549088,0.0010810102355067698,0.0011372628442138308,0.0011867342580300108,0.0012295408339795142,0.0012658227447402998,0.0012957461488201504,0.0013195016209159504,0.0013373001969577845,0.0013493699157382595,0.001355954523788637,0.0013573134214608581,0.0013537200572276192,0.0013454577372516694,0.0013328148472630697,0.0013160876400487337,0.0012955794786071852,0.0012715955672936968,0.0012444355144887226,0.0012144105515198558,0.001181814956554507,0.00114695406560225,0.0011101104561474747,0.0010715828256110285,0.0010316369578531872,9.905471698109832E-4,9.485751242191463E-4,9.059666182415098E-4,8.62955798960464E-4,8.197694451210797E-4,7.766209124107469E-4,7.337077975763362E-4,6.912130516169605E-4,6.493072085284562E-4,6.081483601883429E-4,5.678804755293912E-4,5.286317701011066E-4,4.905157202469902E-4,4.536340834518712E-4,4.180750727639507E-4,3.8391283512202143E-4,3.5120864671016344E-4,3.200137461957706E-4,2.903616395363066E-4,2.6228274935093744E-4,2.3578135519507906E-4,2.108893983098659E-4,1.8755202781569998E-4,1.6580895365819176E-4,1.4561660801765025E-4,1.2693578037493446E-4,1.0973572173158561E-4,9.398288772764757E-5,7.962974039102439E-5,6.662077754901276E-5,5.489773300334159E-5,4.440230106207581E-5,3.5075205134138346E-5,2.685486721875701E-5,1.967652583693631E-5,1.3474034479830275E-5,8.181670695133963E-6,3.7340395101024115E-6,6.773457347335861E-8,-2.8782725794033763E-6,-5.1627963389752305E-6,-6.843685137216114E-6,-7.973763240331752E-6,-8.607316290639185E-6,-8.791028569757087E-6,-9.314227689476197E-5" />
// Retrieval info: 	<generic name="coeffType" value="Signed Binary" />
// Retrieval info: 	<generic name="coeffScaling" value="Auto" />
// Retrieval info: 	<generic name="coeffBitWidth" value="12" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
// Retrieval info: 	<generic name="outType" value="Signed Binary" />
// Retrieval info: 	<generic name="outMSBRound" value="Truncation" />
// Retrieval info: 	<generic name="outMsbBitRem" value="6" />
// Retrieval info: 	<generic name="outLSBRound" value="Truncation" />
// Retrieval info: 	<generic name="outLsbBitRem" value="15" />
// Retrieval info: 	<generic name="resoureEstimation" value="1000,1200,10" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : fir_lpf.vo
// RELATED_FILES: fir_lpf.v, altera_avalon_sc_fifo.v, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, dspba_library_package.vhd, dspba_library.vhd, fir_lpf_0002_rtl.vhd, fir_lpf_0002_ast.vhd, fir_lpf_0002.vhd
